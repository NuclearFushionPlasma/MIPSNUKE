module Ins_MEM(
  input [31:0] Ins_address,
  input clk,reset,
  output[31:0] Ins_output
  );
  assign Ins_output = 0;
endmodule